---------------------------------------------
-- EU Module
--
-- Info:
-- info
--
-- ToDo:
-- ToDo
--
-- Testing:
-- Testing
---------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
---------------------------------------------
entity EU is
    generic(Size : integer := 32);
    port(
        --ToDo
        Clk : in std_logic
    );
end entity EU;
---------------------------------------------
architecture default of EU is
begin
    --ToDo
end default;
---------------------------------------------
