---------------------------------------------
-- FlagRegister Module
--
-- Info:
-- info
--
-- ToDo:
-- ToDo
--
-- Testing:
-- Testing
---------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
---------------------------------------------
entity FlagRegister is
    generic(GenericVariable : integer := GenericValue);
    port(
        --ToDo
    );
end entity FlagRegister;
---------------------------------------------
architecture default of FlagRegister is
begin
    --ToDo
end default;
---------------------------------------------