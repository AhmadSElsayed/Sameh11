---------------------------------------------
-- FlagRegister Module
--
-- Info:
-- info
--
-- ToDo:
-- ToDo
--
-- Testing:
-- Testing
---------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
---------------------------------------------
entity FlagRegister is
    generic(Size : integer := 4);
    port(
        --ToDo
        Clk : in std_logic
    );
end entity FlagRegister;
---------------------------------------------
architecture default of FlagRegister is
begin
    --ToDo
end default;
---------------------------------------------
