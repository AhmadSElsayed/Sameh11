---------------------------------------------
-- CU Module
--
-- Info:
-- info
--
-- ToDo:
-- ToDo
--
-- Testing:
-- Testing
---------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
---------------------------------------------
entity CU is
    port(
        --ToDo
        Clk : in std_logic
    );
end entity CU;
---------------------------------------------
architecture default of CU is
begin
    --ToDo
end default;
---------------------------------------------
