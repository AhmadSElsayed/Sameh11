---------------------------------------------
-- EU Module
--
-- Info:
-- info
--
-- ToDo:
-- ToDo
--
-- Testing:
-- Testing
---------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
---------------------------------------------
entity EU is
    generic(GenericVariable : integer := GenericValue);
    port(
        --ToDo
    );
end entity EU;
---------------------------------------------
architecture default of EU is
begin
    --ToDo
end default;
---------------------------------------------